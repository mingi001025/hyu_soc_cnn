parameter   IN          = 2;  // Number of Input/Output (Batch size)
parameter   ICH         = 3;  // Number of Channel Input 
parameter   OCH         = 2;  // Number of Channel Output

parameter   IX          = 8;  // Number of Input X
parameter   IY          = 4;  // Number of Input Y
parameter	KX			= 4;  // Number of Kernel X
parameter	KY			= 3;  // Number of Kernel Y
parameter   OX          = 5;  // Number of Output X = input X - Kernel X + 1
parameter   OY          = 2;  // Number of Output Y = input Y - kernel Y + 1

parameter	DATA_LEN	= 32; // data length
